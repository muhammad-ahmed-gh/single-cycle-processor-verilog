module immediate_generator (
  
);

endmodule