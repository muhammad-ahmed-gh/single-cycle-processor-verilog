// Instruction Memory, Data Memory & Top-Level Integration
// You will implement:
// A. Instruction Memory
// • Preloaded 
// • Word-aligned addressing
// B. Data Memory
// • Support for ld and sd
// • Word-addressed RAM
// C. CPU Top-Level Module

// You will integrate:
// • PC
// • Instruction memory
// • Control unit
// • Register file
// • ALU
// • Immediate generator
// • Data memory
// • Branch logic
// • All multiplexers and internal wires

// Your responsibilities:
// • Make sure all modules connect correctly
// • Run the full-core simulation
// • Run RISC-V program to test the processor

module data_memory (

);

endmodule