module pc (
  
);

endmodule