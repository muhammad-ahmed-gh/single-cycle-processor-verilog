// Program Counter, Branch Logic & PC Update
// You will design all components related to instruction sequencing:
// • PC register (updates every cycle)
// • PC + 4 adder
// • Branch target calculation
// • Branch decision logic
// • MUX for selecting the next PC
// • Handling branching correctly

// Your responsibilities:
// • Implement PC logic in Verilog
// • Verify correct branching behavior in a testbench

module pc (
  
);

endmodule