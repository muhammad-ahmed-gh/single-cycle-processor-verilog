module top (
  
);

endmodule