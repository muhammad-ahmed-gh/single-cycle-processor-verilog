`timescale 1ns/1ps
module test_bench;
  initial begin

    $display("Hello, world!");

  end
endmodule