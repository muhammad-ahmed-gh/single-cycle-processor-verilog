module test_bench;
  initial begin
    
    $display("Hello, world!");

  end
endmodule