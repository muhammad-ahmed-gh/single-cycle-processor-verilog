// Register File & Immediate Generator
// You will implement: 
// A. Register File 
// • 32 registers 
// • x0 always 0 
// • two read ports, one write port 
// • synchronous write, asynchronous read 
// B. Immediate Generator 
// • Correct extraction and sign-extension of immediates for 
// addi, andi, xori, ori, ld, sd, beq, shift-immediates 

// Your responsibilities: 
// • Implement both modules in Verilog 
// • Create a testbench to verify register reads/writes and immediate formats 

module register_file (
  
);

endmodule