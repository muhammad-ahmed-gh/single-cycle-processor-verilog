// Control Unit (Main Control + ALU Control Merged)
// You will design and implement the Control Unit, responsible for generating all
// internal control signals, including:
// • RegWrite
// • MemWrite
// • MemRead
// • ALUSrc
// • MemToReg
// • Branch
// • ALUControl (merged inside)

// Your responsibilities:
// • Build the control table for all required instructions
// • Implement instruction decoding logic
// • Generate ALUControl directly from opcode + funct3/funct7
// • Provide a testbench that applies opcodes and checks correct control signals

module control_unit (
  
);

endmodule